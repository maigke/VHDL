component and_2 is
  port (
    a : in  std_logic;
    b : in  std_logic;
    c : out std_logic
  );
end component;
